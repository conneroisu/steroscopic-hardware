module compute_SAD #(
    parameter WIN = 3,
    parameter WIN_SIZE = WIN * WIN,
    parameter DATA_SIZE = 8
)(
    
);